.title Spice Simulation 1-1

.include "models/lm2596_5.lib"
.include "models/led_green.lib"
.include "models/s1a.lib"
.include "models/ss24.lib"

*.OPTION ABSTOL=1e-15.
*.OPTION GMIN=1.0e-12.
*.OPTION ITL1=1e5
*.OPTION RSHUNT=1e12
*.OPTION RELTOL=1e-5
*.OPTION GMINSTEPS=1000
*.OPTION ITL3=100

*** V24v    VIN GND 24 AC 24 0 SIN(0V 34V 60Hz)
*** D1      VIN D1_OUT DI_S1A
V12v    VIN GND 12
C1      VIN GND 680uF
XIC1    VIN PWR_5V IC1_OUT GND GND LM2596_5P0_TRANS
XD2     GND IC1_OUT SS24
L1      IC1_OUT PWR_5V 33uH
C2      PWR_5V GND 220uF

*** V24v    VIN GND 24 AC 24 0 SIN(0V 34V 60Hz)
*** D1      VIN D1_OUT DI_S1A
*** C1      D1_OUT GND 100uF
*** XIC1    D1_OUT PWR_5V IC1_OUT GND GND LM2596_5P0_TRANS
*** XD2     GND IC1_OUT SS24
*** L1      IC1_OUT PWR_5V 150uH
*** C2      PWR_5V GND 100uF

*** SIMULATION Commands ***
.tran 1ms 28ms 0 UIC
.control
run
plot v(VIN), v(PWR_5V), v(IC1_OUT)
.endc

.end
