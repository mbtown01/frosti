.title Spice Simulation 1-1

*.OPTION ABSTOL=1e-15.
*.OPTION GMIN=1.0e-12.
*.OPTION ITL1=1e5
*.OPTION RSHUNT=1e12
*.OPTION RELTOL=1e-5
*.OPTION GMINSTEPS=1000
*.OPTION ITL3=100

*SRC=S1A;DI_S1A;Diodes;Si;  50.0V  1.00A  3.00us   Diodes Inc. Rectifier
.MODEL  DI_S1A D  ( IS=7.31e-018 RS=42.0m BV=50.0 IBV=5.00u
+ CJO=42.4p  M=0.333 N=0.775 TT=4.32u )

V1      VIN GND AC 12 0 SIN(0V 30V 10)
D1      VIN D1_OUT DI_S1A
C1      D1_OUT GND 500uF
R1      D1_OUT GND 1

*** SIMULATION Commands ***
.tran 1ms 250ms 0 UIC
.control
run
plot v(D1_OUT), v(VIN)
.endc

.end
